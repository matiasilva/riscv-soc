`ifdef SYNTHESIS
`define SYSFREQ 50000000
`else
`define SYSFREQ 100_000_000
`endif
