/*
	this module produces the required control signal for the ALU
*/

module alucontrol (
	input clk,
	input rst_n,
	input [2:0] alu_op,
	input []
	output [2:0] control
);

endmodule