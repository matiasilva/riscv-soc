module uart_tx(
   input wire clk,
   input wire rst_n,
   input wire [7:0] data.

   output wire sd
);
