`ifdef SYNTHESIS
   `define SYSFREQ 50000000
`else
   `define SYSFREQ 50000000
`endif
